/**************************************************************************
 * Clock Reset UVM Agent
 * Copyright (C) 2024, RISCY-Lib Contributors
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 **************************************************************************/

interface clk_rst_if #(
  parameter NUMBER_OF_CLKS = 1,
  parameter NUMBER_OF_RSTS = 1
);
  logic [NUMBER_OF_CLKS-1:0] clk;
  logic [NUMBER_OF_RSTS-1:0] rst;
  logic [NUMBER_OF_RSTS-1:0] rst_n;

  assign rst_n = ~rst;

endinterface